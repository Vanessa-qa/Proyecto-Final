//Jonathan Garcia Tovar
//Laura Vanessa Quintero Arreola

module ANDbranch
(
	input wire A, B,
	output wire R
);

    assign R = A & B;
	
endmodule